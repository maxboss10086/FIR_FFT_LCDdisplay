library verilog;
use verilog.vl_types.all;
entity spi_dri_tb is
end spi_dri_tb;
